`default_nettype none
module Btn(
    input clk,
	output wire[15:0] out
);

endmodule