/**
 * Demultiplexor:
 * {a, b} = {in, 0} if sel == 0
 *          {0, in} if sel == 1
 */
`default_nettype none

module DMux(
	input wire in,
	input wire sel,
    output wire a,
	output wire b
);

// your implementation comes here:




endmodule
