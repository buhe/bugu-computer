/**
 * 16-way Or: 
 * out = (in[0] or in[1] or ... or in[15])
 */
`default_nettype none

module Or16Way(
	input [15:0] in,
	output out
);




endmodule
