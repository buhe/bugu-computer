`default_nettype none

module Led(
    input clk,
	input wire load,
    output wire led,
	output wire[15:0] out,
	input wire[15:0] in
);
    wire prev;
    Mux MUX(.a(out[0]),.b(in[0]),.sel(load),.out(prev));
    assign led = prev;
	DFFusr DFF1(.clk(clk),.in(prev),.out(out[0]));

endmodule