`default_nettype none
module Led(
    input clk,
	output wire load,
	output wire[15:0] out,
	input wire[15:0] in
);

endmodule